--    Violet
